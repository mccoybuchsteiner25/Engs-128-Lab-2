----------------------------------------------------------------------------
--  Lab 2: AXI Stream FIFO and DMA
----------------------------------------------------------------------------
--  ENGS 128 Spring 2025
--	Author: Kendall Farnham
----------------------------------------------------------------------------
--	Description: AXI Stream FIFO Controller/Responder Interface 
----------------------------------------------------------------------------
-- Library Declarations
library ieee;
use ieee.std_logic_1164.all;

----------------------------------------------------------------------------
-- Entity definition
entity axis_fifo is
	generic (
		DATA_WIDTH	: integer	:= 32;
		FIFO_DEPTH	: integer	:= 1024;
		AC_DATA_WIDTH : integer := 24
	);
	port (
		-- Ports of Axi Responder Bus Interface S00_AXIS
		s00_axis_aclk     : in std_logic;
		s00_axis_aresetn  : in std_logic;
		s00_axis_tready   : out std_logic;
		s00_axis_tdata	  : in std_logic_vector(DATA_WIDTH-1 downto 0);
		s00_axis_tstrb    : in std_logic_vector((DATA_WIDTH/8)-1 downto 0);
		s00_axis_tlast    : in std_logic;
		s00_axis_tvalid   : in std_logic;

		-- Ports of Axi Controller Bus Interface M00_AXIS
		m00_axis_aclk     : in std_logic;
		m00_axis_aresetn  : in std_logic;
		m00_axis_tvalid   : out std_logic;
		m00_axis_tdata    : out std_logic_vector(DATA_WIDTH-1 downto 0);
		m00_axis_tstrb    : out std_logic_vector((DATA_WIDTH/8)-1 downto 0);
		m00_axis_tlast    : out std_logic;
		m00_axis_tready   : in std_logic
	);
end axis_fifo;

----------------------------------------------------------------------------
-- Architecture Definition 
architecture Behavioral of axis_fifo is
----------------------------------------------------------------------------
-- Signals
----------------------------------------------------------------------------  
signal wr_en_s ,rd_en_s : std_logic := '0';
signal wr_data_s, rd_data_s : std_logic_vector(DATA_WIDTH-1 downto 0);
signal empty_s, full_s : std_logic := '0';


----------------------------------------------------------------------------
-- Component Declarations
----------------------------------------------------------------------------  
component fifo is
    Generic (
		FIFO_DEPTH : integer := FIFO_DEPTH;
        DATA_WIDTH : integer := DATA_WIDTH);
    Port ( 
        clk_i       : in std_logic;
        reset_i     : in std_logic;
        
        -- Write channel
        wr_en_i     : in std_logic;
        wr_data_i   : in std_logic_vector(DATA_WIDTH-1 downto 0);
        
        -- Read channel
        rd_en_i     : in std_logic;
        rd_data_o   : out std_logic_vector(DATA_WIDTH-1 downto 0);
        
        -- Status flags
        empty_o         : out std_logic;
        full_o          : out std_logic);   
end component fifo;

----------------------------------------------------------------------------
begin

----------------------------------------------------------------------------
-- Component Instantiations
----------------------------------------------------------------------------   
fifo_stream : fifo
    port map (
        clk_i => s00_axis_aclk,
        reset_i => not s00_axis_aresetn,
        wr_en_i => wr_en_s,
        wr_data_i => wr_data_s,
        rd_en_i => rd_en_s,
        rd_data_o => rd_data_s,
        empty_o => empty_s,
        full_o => full_s);

------------------------------------------------------------------
-- Logic
----------------------------------------------------------------------------  
rd_en_s <= m00_axis_tready and (not empty_s);
wr_en_s <= s00_axis_tvalid and (not full_s);
wr_data_s <= s00_axis_tdata;
s00_axis_tready <= '0' when s00_axis_aresetn = '0' else not full_s;
m00_axis_tdata <= (others=> '0') when s00_axis_aresetn ='0' else rd_data_s;
m00_axis_tvalid <= '0' when m00_axis_aresetn = '0' else not empty_s;
m00_axis_tstrb <= (others => '1'); -- 1111
m00_axis_tlast <= '0'; -- 0



end Behavioral;
